-- MIL-STD-1553 controllers

  constant CFG_GR1553B_ENABLE     : integer := CONFIG_GR1553B_ENABLE;
  constant CFG_GR1553B_RTEN       : integer := CONFIG_GR1553B_RTEN;
  constant CFG_GR1553B_BCEN       : integer := CONFIG_GR1553B_BCEN;
  constant CFG_GR1553B_BMEN       : integer := CONFIG_GR1553B_BMEN;



package version is
  constant grlib_version : integer := 2017200;
  constant grlib_build : integer := 4194;
end;

-- Spacewire interface
  constant CFG_SPWRTR_ENABLE    : integer := CONFIG_SPWRTR_ENABLE;
  constant CFG_SPWRTR_INPUT     : integer := CONFIG_SPWRTR_INPUT;
  constant CFG_SPWRTR_OUTPUT    : integer := CONFIG_SPWRTR_OUTPUT;
  constant CFG_SPWRTR_RTSAME    : integer := CONFIG_SPWRTR_RTSAME;
  constant CFG_SPWRTR_FIFO      : integer := CONFIG_SPWRTR_FIFO;
  constant CFG_SPWRTR_TECHFIFO  : integer := CONFIG_SPWRTR_TECHFIFO;
  constant CFG_SPWRTR_FT        : integer := CONFIG_SPWRTR_FT;
  constant CFG_SPWRTR_SPWEN     : integer := CONFIG_SPWRTR_SPWEN;
  constant CFG_SPWRTR_AMBAEN    : integer := CONFIG_SPWRTR_AMBAEN;
  constant CFG_SPWRTR_FIFOEN    : integer := CONFIG_SPWRTR_FIFOEN;
  constant CFG_SPWRTR_SPWPORTS  : integer := CONFIG_SPWRTR_SPWPORTS;
  constant CFG_SPWRTR_AMBAPORTS : integer := CONFIG_SPWRTR_AMBAPORTS;
  constant CFG_SPWRTR_FIFOPORTS : integer := CONFIG_SPWRTR_FIFOPORTS;
  constant CFG_SPWRTR_ARB       : integer := CONFIG_SPWRTR_ARB;
  constant CFG_SPWRTR_RMAP      : integer := CONFIG_SPWRTR_RMAP;
  constant CFG_SPWRTR_RMAPCRC   : integer := CONFIG_SPWRTR_RMAPCRC;
  constant CFG_SPWRTR_FIFO2     : integer := CONFIG_SPWRTR_FIFO2;
  constant CFG_SPWRTR_ALMOST    : integer := CONFIG_SPWRTR_ALMOST;
  constant CFG_SPWRTR_RXUNAL    : integer := CONFIG_SPWRTR_RXUNAL;
  constant CFG_SPWRTR_RMAPBUF   : integer := CONFIG_SPWRTR_RMAPBUF;
  constant CFG_SPWRTR_DMACHAN   : integer := CONFIG_SPWRTR_DMACHAN;
  constant CFG_SPWRTR_AHBSLVEN  : integer := CONFIG_SPWRTR_AHBSLVEN;
  constant CFG_SPWRTR_TIMERBITS : integer := CONFIG_SPWRTR_TIMERBITS;
  constant CFG_SPWRTR_PNP       : integer := CONFIG_SPWRTR_PNP;
  constant CFG_SPWRTR_AUTOSCRUB : integer := CONFIG_SPWRTR_AUTOSCRUB;


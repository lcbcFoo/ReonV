-- Dynamic Partial Reconfiguration
  constant CFG_PRC : integer := CONFIG_PARTIAL;
  constant CFG_CRC_EN : integer := CONFIG_CRC;
  constant CFG_EDAC_EN : integer := CONFIG_EDAC;
  constant CFG_WORDS_BLOCK : integer := CONFIG_BLOCK;
  constant CFG_DCM_FIFO : integer := CONFIG_DCM_FIFO;
  constant CFG_DPR_FIFO : integer := CFG_DPRFIFO;


package vcomponents is
end;

